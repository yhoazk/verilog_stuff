module fsm_0
